import Vector::*;
import Pipe::*;
import MemTypes::*;
import ConnectalConfig::*;
import DmaConfig::*;

`include "ConnectalProjectConfig.bsv"
typedef `NumChannels NumChannels;

interface DmaTopPins;
   // derived from pcie clock
   interface Clock clock;
   interface Reset reset;
   // data out to application logic
   interface Vector#(NumChannels,PipeOut#(MemDataF#(DataBusWidth))) readData;
   // data in from application logic
   interface Vector#(NumChannels,PipeIn#(MemDataF#(DataBusWidth)))  writeData;
endinterface
